module frownyFace_tb();

logic [15:0][15:0]Grn;
frownyFace dut(.*);
initial begin 




#10;

$stop;


end



endmodule 