module test(
);

always_comb begin 
	dsfsf
	dsfsf

	case(balls) 


		dsfsf
	endcase
	
	
end