module frownyFace(

output logic [15:0][15:0]Grn
);


always_comb begin

	 Grn[0] = 16'b1111111111111111;	
	 Grn[1] = 16'b1000000000000001;
	 Grn[2] = 16'b1000000000001101;	
	 Grn[3] = 16'b1001110000111001;
	 Grn[4] = 16'b1001010000100001;		
	 Grn[5] = 16'b1001110000100001;		
	 Grn[6] = 16'b1000000000100001;		
	 Grn[7] = 16'b1000000000100001;		
	 Grn[8] = 16'b1000000000100001;		
	 Grn[9] = 16'b1000000000100001;		
	Grn[10] = 16'b1001110000100001;		
	Grn[11] = 16'b1001010000100001;		
	Grn[12] = 16'b1001110000111001;		
	Grn[13] = 16'b1000000000001101;		
	Grn[14] = 16'b1000000000000001;		
	Grn[15] = 16'b1111111111111111;		


	end










endmodule 
